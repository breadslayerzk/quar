library verilog;
use verilog.vl_types.all;
entity complee_vlg_vec_tst is
end complee_vlg_vec_tst;
