library verilog;
use verilog.vl_types.all;
entity comple_vlg_vec_tst is
end comple_vlg_vec_tst;
